<svg width="24" height="24" viewBox="0 0 24 24" fill="none" xmlns="http://www.w3.org/2000/svg">
<path d="M11.9999 2.40002C9.5999 2.40002 7.9999 3.20002 7.9999 3.20002C7.9999 3.20002 7.1999 4.80002 7.1999 8.00002H7.2999C7.4247 8.54882 7.62178 8.9719 7.62178 8.9719C7.45218 9.0695 7.17325 9.37931 7.24365 9.92971C7.37485 10.9561 7.81983 11.2159 8.10303 11.2375C8.21103 12.1959 9.2399 13.4216 9.5999 13.6V15.2C9.59815 15.2053 9.5939 15.2089 9.59209 15.2141C9.32753 15.2469 9.0915 15.403 8.97178 15.6453L8.72178 16.1485C6.74734 17.2556 2.3999 16.9811 2.3999 21.6H21.5999C21.5999 16.9811 17.2525 17.2556 15.278 16.1485L15.028 15.6453C14.9083 15.403 14.6723 15.2469 14.4077 15.2141C14.4059 15.2089 14.4017 15.2053 14.3999 15.2V13.6C14.7599 13.4216 15.7888 12.1967 15.8968 11.2391C16.18 11.2175 16.625 10.9561 16.7562 9.92971C16.8266 9.37851 16.5476 9.0695 16.378 8.9719L16.7077 8.00002H16.7999C16.7999 5.60002 15.9999 3.20002 15.9999 3.20002C15.9999 3.20002 14.3999 2.40002 11.9999 2.40002ZM11.9999 3.20002C12.4415 3.20002 12.7999 3.55842 12.7999 4.00002V4.80002H13.5999C14.0415 4.80002 14.3999 5.15842 14.3999 5.60002C14.3999 6.04162 14.0415 6.40002 13.5999 6.40002H12.7999V7.20002C12.7999 7.64162 12.4415 8.00002 11.9999 8.00002C11.5583 8.00002 11.1999 7.64162 11.1999 7.20002V6.40002H10.3999C9.9583 6.40002 9.5999 6.04162 9.5999 5.60002C9.5999 5.15842 9.9583 4.80002 10.3999 4.80002H11.1999V4.00002C11.1999 3.55842 11.5583 3.20002 11.9999 3.20002Z" fill="white"/>
</svg>